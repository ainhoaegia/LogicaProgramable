-- PROYECTO LÓGICA PROGRAMABLE
